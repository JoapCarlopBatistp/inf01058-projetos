library verilog;
use verilog.vl_types.all;
entity Trabalho_Final_vlg_vec_tst is
end Trabalho_Final_vlg_vec_tst;
